module Clmul(
  input  [31:0] io_A_in,
  input  [31:0] io_B_in,
  output [31:0] io_C_out
);
  wire [31:0] terms_0 = io_B_in[0] ? io_A_in : 32'h0; // @[ZbcExt.scala 19:8]
  wire [32:0] terms_shifted_1 = {io_A_in, 1'h0}; // @[ZbcExt.scala 18:28]
  wire [32:0] terms_1 = io_B_in[1] ? terms_shifted_1 : 33'h0; // @[ZbcExt.scala 19:8]
  wire [33:0] terms_shifted_2 = {io_A_in, 2'h0}; // @[ZbcExt.scala 18:28]
  wire [33:0] terms_2 = io_B_in[2] ? terms_shifted_2 : 34'h0; // @[ZbcExt.scala 19:8]
  wire [34:0] terms_shifted_3 = {io_A_in, 3'h0}; // @[ZbcExt.scala 18:28]
  wire [34:0] terms_3 = io_B_in[3] ? terms_shifted_3 : 35'h0; // @[ZbcExt.scala 19:8]
  wire [35:0] terms_shifted_4 = {io_A_in, 4'h0}; // @[ZbcExt.scala 18:28]
  wire [35:0] terms_4 = io_B_in[4] ? terms_shifted_4 : 36'h0; // @[ZbcExt.scala 19:8]
  wire [36:0] terms_shifted_5 = {io_A_in, 5'h0}; // @[ZbcExt.scala 18:28]
  wire [36:0] terms_5 = io_B_in[5] ? terms_shifted_5 : 37'h0; // @[ZbcExt.scala 19:8]
  wire [37:0] terms_shifted_6 = {io_A_in, 6'h0}; // @[ZbcExt.scala 18:28]
  wire [37:0] terms_6 = io_B_in[6] ? terms_shifted_6 : 38'h0; // @[ZbcExt.scala 19:8]
  wire [38:0] terms_shifted_7 = {io_A_in, 7'h0}; // @[ZbcExt.scala 18:28]
  wire [38:0] terms_7 = io_B_in[7] ? terms_shifted_7 : 39'h0; // @[ZbcExt.scala 19:8]
  wire [39:0] terms_shifted_8 = {io_A_in, 8'h0}; // @[ZbcExt.scala 18:28]
  wire [39:0] terms_8 = io_B_in[8] ? terms_shifted_8 : 40'h0; // @[ZbcExt.scala 19:8]
  wire [40:0] terms_shifted_9 = {io_A_in, 9'h0}; // @[ZbcExt.scala 18:28]
  wire [40:0] terms_9 = io_B_in[9] ? terms_shifted_9 : 41'h0; // @[ZbcExt.scala 19:8]
  wire [41:0] terms_shifted_10 = {io_A_in, 10'h0}; // @[ZbcExt.scala 18:28]
  wire [41:0] terms_10 = io_B_in[10] ? terms_shifted_10 : 42'h0; // @[ZbcExt.scala 19:8]
  wire [42:0] terms_shifted_11 = {io_A_in, 11'h0}; // @[ZbcExt.scala 18:28]
  wire [42:0] terms_11 = io_B_in[11] ? terms_shifted_11 : 43'h0; // @[ZbcExt.scala 19:8]
  wire [43:0] terms_shifted_12 = {io_A_in, 12'h0}; // @[ZbcExt.scala 18:28]
  wire [43:0] terms_12 = io_B_in[12] ? terms_shifted_12 : 44'h0; // @[ZbcExt.scala 19:8]
  wire [44:0] terms_shifted_13 = {io_A_in, 13'h0}; // @[ZbcExt.scala 18:28]
  wire [44:0] terms_13 = io_B_in[13] ? terms_shifted_13 : 45'h0; // @[ZbcExt.scala 19:8]
  wire [45:0] terms_shifted_14 = {io_A_in, 14'h0}; // @[ZbcExt.scala 18:28]
  wire [45:0] terms_14 = io_B_in[14] ? terms_shifted_14 : 46'h0; // @[ZbcExt.scala 19:8]
  wire [46:0] terms_shifted_15 = {io_A_in, 15'h0}; // @[ZbcExt.scala 18:28]
  wire [46:0] terms_15 = io_B_in[15] ? terms_shifted_15 : 47'h0; // @[ZbcExt.scala 19:8]
  wire [47:0] terms_shifted_16 = {io_A_in, 16'h0}; // @[ZbcExt.scala 18:28]
  wire [47:0] terms_16 = io_B_in[16] ? terms_shifted_16 : 48'h0; // @[ZbcExt.scala 19:8]
  wire [48:0] terms_shifted_17 = {io_A_in, 17'h0}; // @[ZbcExt.scala 18:28]
  wire [48:0] terms_17 = io_B_in[17] ? terms_shifted_17 : 49'h0; // @[ZbcExt.scala 19:8]
  wire [49:0] terms_shifted_18 = {io_A_in, 18'h0}; // @[ZbcExt.scala 18:28]
  wire [49:0] terms_18 = io_B_in[18] ? terms_shifted_18 : 50'h0; // @[ZbcExt.scala 19:8]
  wire [50:0] terms_shifted_19 = {io_A_in, 19'h0}; // @[ZbcExt.scala 18:28]
  wire [50:0] terms_19 = io_B_in[19] ? terms_shifted_19 : 51'h0; // @[ZbcExt.scala 19:8]
  wire [51:0] terms_shifted_20 = {io_A_in, 20'h0}; // @[ZbcExt.scala 18:28]
  wire [51:0] terms_20 = io_B_in[20] ? terms_shifted_20 : 52'h0; // @[ZbcExt.scala 19:8]
  wire [52:0] terms_shifted_21 = {io_A_in, 21'h0}; // @[ZbcExt.scala 18:28]
  wire [52:0] terms_21 = io_B_in[21] ? terms_shifted_21 : 53'h0; // @[ZbcExt.scala 19:8]
  wire [53:0] terms_shifted_22 = {io_A_in, 22'h0}; // @[ZbcExt.scala 18:28]
  wire [53:0] terms_22 = io_B_in[22] ? terms_shifted_22 : 54'h0; // @[ZbcExt.scala 19:8]
  wire [54:0] terms_shifted_23 = {io_A_in, 23'h0}; // @[ZbcExt.scala 18:28]
  wire [54:0] terms_23 = io_B_in[23] ? terms_shifted_23 : 55'h0; // @[ZbcExt.scala 19:8]
  wire [55:0] terms_shifted_24 = {io_A_in, 24'h0}; // @[ZbcExt.scala 18:28]
  wire [55:0] terms_24 = io_B_in[24] ? terms_shifted_24 : 56'h0; // @[ZbcExt.scala 19:8]
  wire [56:0] terms_shifted_25 = {io_A_in, 25'h0}; // @[ZbcExt.scala 18:28]
  wire [56:0] terms_25 = io_B_in[25] ? terms_shifted_25 : 57'h0; // @[ZbcExt.scala 19:8]
  wire [57:0] terms_shifted_26 = {io_A_in, 26'h0}; // @[ZbcExt.scala 18:28]
  wire [57:0] terms_26 = io_B_in[26] ? terms_shifted_26 : 58'h0; // @[ZbcExt.scala 19:8]
  wire [58:0] terms_shifted_27 = {io_A_in, 27'h0}; // @[ZbcExt.scala 18:28]
  wire [58:0] terms_27 = io_B_in[27] ? terms_shifted_27 : 59'h0; // @[ZbcExt.scala 19:8]
  wire [59:0] terms_shifted_28 = {io_A_in, 28'h0}; // @[ZbcExt.scala 18:28]
  wire [59:0] terms_28 = io_B_in[28] ? terms_shifted_28 : 60'h0; // @[ZbcExt.scala 19:8]
  wire [60:0] terms_shifted_29 = {io_A_in, 29'h0}; // @[ZbcExt.scala 18:28]
  wire [60:0] terms_29 = io_B_in[29] ? terms_shifted_29 : 61'h0; // @[ZbcExt.scala 19:8]
  wire [61:0] terms_shifted_30 = {io_A_in, 30'h0}; // @[ZbcExt.scala 18:28]
  wire [61:0] terms_30 = io_B_in[30] ? terms_shifted_30 : 62'h0; // @[ZbcExt.scala 19:8]
  wire [32:0] _GEN_0 = {{1'd0}, terms_0}; // @[ZbcExt.scala 23:30]
  wire [32:0] _io_C_out_T = _GEN_0 ^ terms_1; // @[ZbcExt.scala 23:30]
  wire [33:0] _GEN_1 = {{1'd0}, _io_C_out_T}; // @[ZbcExt.scala 23:30]
  wire [33:0] _io_C_out_T_1 = _GEN_1 ^ terms_2; // @[ZbcExt.scala 23:30]
  wire [34:0] _GEN_2 = {{1'd0}, _io_C_out_T_1}; // @[ZbcExt.scala 23:30]
  wire [34:0] _io_C_out_T_2 = _GEN_2 ^ terms_3; // @[ZbcExt.scala 23:30]
  wire [35:0] _GEN_3 = {{1'd0}, _io_C_out_T_2}; // @[ZbcExt.scala 23:30]
  wire [35:0] _io_C_out_T_3 = _GEN_3 ^ terms_4; // @[ZbcExt.scala 23:30]
  wire [36:0] _GEN_4 = {{1'd0}, _io_C_out_T_3}; // @[ZbcExt.scala 23:30]
  wire [36:0] _io_C_out_T_4 = _GEN_4 ^ terms_5; // @[ZbcExt.scala 23:30]
  wire [37:0] _GEN_5 = {{1'd0}, _io_C_out_T_4}; // @[ZbcExt.scala 23:30]
  wire [37:0] _io_C_out_T_5 = _GEN_5 ^ terms_6; // @[ZbcExt.scala 23:30]
  wire [38:0] _GEN_6 = {{1'd0}, _io_C_out_T_5}; // @[ZbcExt.scala 23:30]
  wire [38:0] _io_C_out_T_6 = _GEN_6 ^ terms_7; // @[ZbcExt.scala 23:30]
  wire [39:0] _GEN_7 = {{1'd0}, _io_C_out_T_6}; // @[ZbcExt.scala 23:30]
  wire [39:0] _io_C_out_T_7 = _GEN_7 ^ terms_8; // @[ZbcExt.scala 23:30]
  wire [40:0] _GEN_8 = {{1'd0}, _io_C_out_T_7}; // @[ZbcExt.scala 23:30]
  wire [40:0] _io_C_out_T_8 = _GEN_8 ^ terms_9; // @[ZbcExt.scala 23:30]
  wire [41:0] _GEN_9 = {{1'd0}, _io_C_out_T_8}; // @[ZbcExt.scala 23:30]
  wire [41:0] _io_C_out_T_9 = _GEN_9 ^ terms_10; // @[ZbcExt.scala 23:30]
  wire [42:0] _GEN_10 = {{1'd0}, _io_C_out_T_9}; // @[ZbcExt.scala 23:30]
  wire [42:0] _io_C_out_T_10 = _GEN_10 ^ terms_11; // @[ZbcExt.scala 23:30]
  wire [43:0] _GEN_11 = {{1'd0}, _io_C_out_T_10}; // @[ZbcExt.scala 23:30]
  wire [43:0] _io_C_out_T_11 = _GEN_11 ^ terms_12; // @[ZbcExt.scala 23:30]
  wire [44:0] _GEN_12 = {{1'd0}, _io_C_out_T_11}; // @[ZbcExt.scala 23:30]
  wire [44:0] _io_C_out_T_12 = _GEN_12 ^ terms_13; // @[ZbcExt.scala 23:30]
  wire [45:0] _GEN_13 = {{1'd0}, _io_C_out_T_12}; // @[ZbcExt.scala 23:30]
  wire [45:0] _io_C_out_T_13 = _GEN_13 ^ terms_14; // @[ZbcExt.scala 23:30]
  wire [46:0] _GEN_14 = {{1'd0}, _io_C_out_T_13}; // @[ZbcExt.scala 23:30]
  wire [46:0] _io_C_out_T_14 = _GEN_14 ^ terms_15; // @[ZbcExt.scala 23:30]
  wire [47:0] _GEN_15 = {{1'd0}, _io_C_out_T_14}; // @[ZbcExt.scala 23:30]
  wire [47:0] _io_C_out_T_15 = _GEN_15 ^ terms_16; // @[ZbcExt.scala 23:30]
  wire [48:0] _GEN_16 = {{1'd0}, _io_C_out_T_15}; // @[ZbcExt.scala 23:30]
  wire [48:0] _io_C_out_T_16 = _GEN_16 ^ terms_17; // @[ZbcExt.scala 23:30]
  wire [49:0] _GEN_17 = {{1'd0}, _io_C_out_T_16}; // @[ZbcExt.scala 23:30]
  wire [49:0] _io_C_out_T_17 = _GEN_17 ^ terms_18; // @[ZbcExt.scala 23:30]
  wire [50:0] _GEN_18 = {{1'd0}, _io_C_out_T_17}; // @[ZbcExt.scala 23:30]
  wire [50:0] _io_C_out_T_18 = _GEN_18 ^ terms_19; // @[ZbcExt.scala 23:30]
  wire [51:0] _GEN_19 = {{1'd0}, _io_C_out_T_18}; // @[ZbcExt.scala 23:30]
  wire [51:0] _io_C_out_T_19 = _GEN_19 ^ terms_20; // @[ZbcExt.scala 23:30]
  wire [52:0] _GEN_20 = {{1'd0}, _io_C_out_T_19}; // @[ZbcExt.scala 23:30]
  wire [52:0] _io_C_out_T_20 = _GEN_20 ^ terms_21; // @[ZbcExt.scala 23:30]
  wire [53:0] _GEN_21 = {{1'd0}, _io_C_out_T_20}; // @[ZbcExt.scala 23:30]
  wire [53:0] _io_C_out_T_21 = _GEN_21 ^ terms_22; // @[ZbcExt.scala 23:30]
  wire [54:0] _GEN_22 = {{1'd0}, _io_C_out_T_21}; // @[ZbcExt.scala 23:30]
  wire [54:0] _io_C_out_T_22 = _GEN_22 ^ terms_23; // @[ZbcExt.scala 23:30]
  wire [55:0] _GEN_23 = {{1'd0}, _io_C_out_T_22}; // @[ZbcExt.scala 23:30]
  wire [55:0] _io_C_out_T_23 = _GEN_23 ^ terms_24; // @[ZbcExt.scala 23:30]
  wire [56:0] _GEN_24 = {{1'd0}, _io_C_out_T_23}; // @[ZbcExt.scala 23:30]
  wire [56:0] _io_C_out_T_24 = _GEN_24 ^ terms_25; // @[ZbcExt.scala 23:30]
  wire [57:0] _GEN_25 = {{1'd0}, _io_C_out_T_24}; // @[ZbcExt.scala 23:30]
  wire [57:0] _io_C_out_T_25 = _GEN_25 ^ terms_26; // @[ZbcExt.scala 23:30]
  wire [58:0] _GEN_26 = {{1'd0}, _io_C_out_T_25}; // @[ZbcExt.scala 23:30]
  wire [58:0] _io_C_out_T_26 = _GEN_26 ^ terms_27; // @[ZbcExt.scala 23:30]
  wire [59:0] _GEN_27 = {{1'd0}, _io_C_out_T_26}; // @[ZbcExt.scala 23:30]
  wire [59:0] _io_C_out_T_27 = _GEN_27 ^ terms_28; // @[ZbcExt.scala 23:30]
  wire [60:0] _GEN_28 = {{1'd0}, _io_C_out_T_27}; // @[ZbcExt.scala 23:30]
  wire [60:0] _io_C_out_T_28 = _GEN_28 ^ terms_29; // @[ZbcExt.scala 23:30]
  wire [61:0] _GEN_29 = {{1'd0}, _io_C_out_T_28}; // @[ZbcExt.scala 23:30]
  wire [61:0] _io_C_out_T_29 = _GEN_29 ^ terms_30; // @[ZbcExt.scala 23:30]
  assign io_C_out = _io_C_out_T_29[31:0]; // @[ZbcExt.scala 23:12]
endmodule
module Clmulh(
  input  [31:0] io_A_in,
  input  [31:0] io_B_in,
  output [31:0] io_C_out
);
  wire [31:0] terms_shifted = {{31'd0}, io_A_in[31]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_0 = io_B_in[1] ? terms_shifted : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_1 = {{30'd0}, io_A_in[31:30]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_1 = io_B_in[2] ? terms_shifted_1 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_2 = {{29'd0}, io_A_in[31:29]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_2 = io_B_in[3] ? terms_shifted_2 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_3 = {{28'd0}, io_A_in[31:28]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_3 = io_B_in[4] ? terms_shifted_3 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_4 = {{27'd0}, io_A_in[31:27]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_4 = io_B_in[5] ? terms_shifted_4 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_5 = {{26'd0}, io_A_in[31:26]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_5 = io_B_in[6] ? terms_shifted_5 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_6 = {{25'd0}, io_A_in[31:25]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_6 = io_B_in[7] ? terms_shifted_6 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_7 = {{24'd0}, io_A_in[31:24]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_7 = io_B_in[8] ? terms_shifted_7 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_8 = {{23'd0}, io_A_in[31:23]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_8 = io_B_in[9] ? terms_shifted_8 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_9 = {{22'd0}, io_A_in[31:22]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_9 = io_B_in[10] ? terms_shifted_9 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_10 = {{21'd0}, io_A_in[31:21]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_10 = io_B_in[11] ? terms_shifted_10 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_11 = {{20'd0}, io_A_in[31:20]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_11 = io_B_in[12] ? terms_shifted_11 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_12 = {{19'd0}, io_A_in[31:19]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_12 = io_B_in[13] ? terms_shifted_12 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_13 = {{18'd0}, io_A_in[31:18]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_13 = io_B_in[14] ? terms_shifted_13 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_14 = {{17'd0}, io_A_in[31:17]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_14 = io_B_in[15] ? terms_shifted_14 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_15 = {{16'd0}, io_A_in[31:16]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_15 = io_B_in[16] ? terms_shifted_15 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_16 = {{15'd0}, io_A_in[31:15]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_16 = io_B_in[17] ? terms_shifted_16 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_17 = {{14'd0}, io_A_in[31:14]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_17 = io_B_in[18] ? terms_shifted_17 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_18 = {{13'd0}, io_A_in[31:13]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_18 = io_B_in[19] ? terms_shifted_18 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_19 = {{12'd0}, io_A_in[31:12]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_19 = io_B_in[20] ? terms_shifted_19 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_20 = {{11'd0}, io_A_in[31:11]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_20 = io_B_in[21] ? terms_shifted_20 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_21 = {{10'd0}, io_A_in[31:10]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_21 = io_B_in[22] ? terms_shifted_21 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_22 = {{9'd0}, io_A_in[31:9]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_22 = io_B_in[23] ? terms_shifted_22 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_23 = {{8'd0}, io_A_in[31:8]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_23 = io_B_in[24] ? terms_shifted_23 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_24 = {{7'd0}, io_A_in[31:7]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_24 = io_B_in[25] ? terms_shifted_24 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_25 = {{6'd0}, io_A_in[31:6]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_25 = io_B_in[26] ? terms_shifted_25 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_26 = {{5'd0}, io_A_in[31:5]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_26 = io_B_in[27] ? terms_shifted_26 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_27 = {{4'd0}, io_A_in[31:4]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_27 = io_B_in[28] ? terms_shifted_27 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_28 = {{3'd0}, io_A_in[31:3]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_28 = io_B_in[29] ? terms_shifted_28 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_29 = {{2'd0}, io_A_in[31:2]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_29 = io_B_in[30] ? terms_shifted_29 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] terms_shifted_30 = {{1'd0}, io_A_in[31:1]}; // @[ZbcExt.scala 36:27]
  wire [31:0] terms_30 = io_B_in[31] ? terms_shifted_30 : 32'h0; // @[ZbcExt.scala 37:8]
  wire [31:0] _io_C_out_T = terms_0 ^ terms_1; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_1 = _io_C_out_T ^ terms_2; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_2 = _io_C_out_T_1 ^ terms_3; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_3 = _io_C_out_T_2 ^ terms_4; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_4 = _io_C_out_T_3 ^ terms_5; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_5 = _io_C_out_T_4 ^ terms_6; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_6 = _io_C_out_T_5 ^ terms_7; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_7 = _io_C_out_T_6 ^ terms_8; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_8 = _io_C_out_T_7 ^ terms_9; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_9 = _io_C_out_T_8 ^ terms_10; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_10 = _io_C_out_T_9 ^ terms_11; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_11 = _io_C_out_T_10 ^ terms_12; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_12 = _io_C_out_T_11 ^ terms_13; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_13 = _io_C_out_T_12 ^ terms_14; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_14 = _io_C_out_T_13 ^ terms_15; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_15 = _io_C_out_T_14 ^ terms_16; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_16 = _io_C_out_T_15 ^ terms_17; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_17 = _io_C_out_T_16 ^ terms_18; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_18 = _io_C_out_T_17 ^ terms_19; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_19 = _io_C_out_T_18 ^ terms_20; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_20 = _io_C_out_T_19 ^ terms_21; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_21 = _io_C_out_T_20 ^ terms_22; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_22 = _io_C_out_T_21 ^ terms_23; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_23 = _io_C_out_T_22 ^ terms_24; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_24 = _io_C_out_T_23 ^ terms_25; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_25 = _io_C_out_T_24 ^ terms_26; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_26 = _io_C_out_T_25 ^ terms_27; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_27 = _io_C_out_T_26 ^ terms_28; // @[ZbcExt.scala 41:30]
  wire [31:0] _io_C_out_T_28 = _io_C_out_T_27 ^ terms_29; // @[ZbcExt.scala 41:30]
  assign io_C_out = _io_C_out_T_28 ^ terms_30; // @[ZbcExt.scala 41:30]
endmodule
module Clmulr(
  input  [31:0] io_A_in,
  input  [31:0] io_B_in,
  output [31:0] io_C_out
);
  wire [31:0] terms_shifted = {{31'd0}, io_A_in[31]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_0 = io_B_in[0] ? terms_shifted : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_1 = {{30'd0}, io_A_in[31:30]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_1 = io_B_in[1] ? terms_shifted_1 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_2 = {{29'd0}, io_A_in[31:29]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_2 = io_B_in[2] ? terms_shifted_2 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_3 = {{28'd0}, io_A_in[31:28]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_3 = io_B_in[3] ? terms_shifted_3 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_4 = {{27'd0}, io_A_in[31:27]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_4 = io_B_in[4] ? terms_shifted_4 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_5 = {{26'd0}, io_A_in[31:26]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_5 = io_B_in[5] ? terms_shifted_5 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_6 = {{25'd0}, io_A_in[31:25]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_6 = io_B_in[6] ? terms_shifted_6 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_7 = {{24'd0}, io_A_in[31:24]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_7 = io_B_in[7] ? terms_shifted_7 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_8 = {{23'd0}, io_A_in[31:23]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_8 = io_B_in[8] ? terms_shifted_8 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_9 = {{22'd0}, io_A_in[31:22]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_9 = io_B_in[9] ? terms_shifted_9 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_10 = {{21'd0}, io_A_in[31:21]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_10 = io_B_in[10] ? terms_shifted_10 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_11 = {{20'd0}, io_A_in[31:20]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_11 = io_B_in[11] ? terms_shifted_11 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_12 = {{19'd0}, io_A_in[31:19]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_12 = io_B_in[12] ? terms_shifted_12 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_13 = {{18'd0}, io_A_in[31:18]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_13 = io_B_in[13] ? terms_shifted_13 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_14 = {{17'd0}, io_A_in[31:17]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_14 = io_B_in[14] ? terms_shifted_14 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_15 = {{16'd0}, io_A_in[31:16]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_15 = io_B_in[15] ? terms_shifted_15 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_16 = {{15'd0}, io_A_in[31:15]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_16 = io_B_in[16] ? terms_shifted_16 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_17 = {{14'd0}, io_A_in[31:14]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_17 = io_B_in[17] ? terms_shifted_17 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_18 = {{13'd0}, io_A_in[31:13]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_18 = io_B_in[18] ? terms_shifted_18 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_19 = {{12'd0}, io_A_in[31:12]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_19 = io_B_in[19] ? terms_shifted_19 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_20 = {{11'd0}, io_A_in[31:11]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_20 = io_B_in[20] ? terms_shifted_20 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_21 = {{10'd0}, io_A_in[31:10]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_21 = io_B_in[21] ? terms_shifted_21 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_22 = {{9'd0}, io_A_in[31:9]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_22 = io_B_in[22] ? terms_shifted_22 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_23 = {{8'd0}, io_A_in[31:8]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_23 = io_B_in[23] ? terms_shifted_23 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_24 = {{7'd0}, io_A_in[31:7]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_24 = io_B_in[24] ? terms_shifted_24 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_25 = {{6'd0}, io_A_in[31:6]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_25 = io_B_in[25] ? terms_shifted_25 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_26 = {{5'd0}, io_A_in[31:5]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_26 = io_B_in[26] ? terms_shifted_26 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_27 = {{4'd0}, io_A_in[31:4]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_27 = io_B_in[27] ? terms_shifted_27 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_28 = {{3'd0}, io_A_in[31:3]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_28 = io_B_in[28] ? terms_shifted_28 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_29 = {{2'd0}, io_A_in[31:2]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_29 = io_B_in[29] ? terms_shifted_29 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] terms_shifted_30 = {{1'd0}, io_A_in[31:1]}; // @[ZbcExt.scala 56:27]
  wire [31:0] terms_30 = io_B_in[30] ? terms_shifted_30 : 32'h0; // @[ZbcExt.scala 57:8]
  wire [31:0] _io_C_out_T = terms_0 ^ terms_1; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_1 = _io_C_out_T ^ terms_2; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_2 = _io_C_out_T_1 ^ terms_3; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_3 = _io_C_out_T_2 ^ terms_4; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_4 = _io_C_out_T_3 ^ terms_5; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_5 = _io_C_out_T_4 ^ terms_6; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_6 = _io_C_out_T_5 ^ terms_7; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_7 = _io_C_out_T_6 ^ terms_8; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_8 = _io_C_out_T_7 ^ terms_9; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_9 = _io_C_out_T_8 ^ terms_10; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_10 = _io_C_out_T_9 ^ terms_11; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_11 = _io_C_out_T_10 ^ terms_12; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_12 = _io_C_out_T_11 ^ terms_13; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_13 = _io_C_out_T_12 ^ terms_14; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_14 = _io_C_out_T_13 ^ terms_15; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_15 = _io_C_out_T_14 ^ terms_16; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_16 = _io_C_out_T_15 ^ terms_17; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_17 = _io_C_out_T_16 ^ terms_18; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_18 = _io_C_out_T_17 ^ terms_19; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_19 = _io_C_out_T_18 ^ terms_20; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_20 = _io_C_out_T_19 ^ terms_21; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_21 = _io_C_out_T_20 ^ terms_22; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_22 = _io_C_out_T_21 ^ terms_23; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_23 = _io_C_out_T_22 ^ terms_24; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_24 = _io_C_out_T_23 ^ terms_25; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_25 = _io_C_out_T_24 ^ terms_26; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_26 = _io_C_out_T_25 ^ terms_27; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_27 = _io_C_out_T_26 ^ terms_28; // @[ZbcExt.scala 61:30]
  wire [31:0] _io_C_out_T_28 = _io_C_out_T_27 ^ terms_29; // @[ZbcExt.scala 61:30]
  assign io_C_out = _io_C_out_T_28 ^ terms_30; // @[ZbcExt.scala 61:30]
endmodule
module Zbc(
  input         clock,
  input         reset,
  input  [31:0] io_rs1,
  input  [31:0] io_rs2,
  input  [1:0]  io_INSTR_SEL,
  output [31:0] io_rd
);
  wire [31:0] CLMUL_io_A_in; // @[ZbcExt.scala 75:21]
  wire [31:0] CLMUL_io_B_in; // @[ZbcExt.scala 75:21]
  wire [31:0] CLMUL_io_C_out; // @[ZbcExt.scala 75:21]
  wire [31:0] CLMULH_io_A_in; // @[ZbcExt.scala 77:22]
  wire [31:0] CLMULH_io_B_in; // @[ZbcExt.scala 77:22]
  wire [31:0] CLMULH_io_C_out; // @[ZbcExt.scala 77:22]
  wire [31:0] CLMULR_io_A_in; // @[ZbcExt.scala 79:22]
  wire [31:0] CLMULR_io_B_in; // @[ZbcExt.scala 79:22]
  wire [31:0] CLMULR_io_C_out; // @[ZbcExt.scala 79:22]
  wire [31:0] _GEN_0 = 2'h2 == io_INSTR_SEL ? io_rs1 : 32'h0; // @[ZbcExt.scala 104:22 87:18 92:24]
  wire [31:0] _GEN_1 = 2'h2 == io_INSTR_SEL ? io_rs2 : 32'h0; // @[ZbcExt.scala 105:22 88:18 92:24]
  wire [31:0] _GEN_2 = 2'h2 == io_INSTR_SEL ? CLMULR_io_C_out : 32'h0; // @[ZbcExt.scala 106:10 92:24]
  wire [31:0] _GEN_3 = 2'h1 == io_INSTR_SEL ? io_rs1 : 32'h0; // @[ZbcExt.scala 84:18 92:24 99:22]
  wire [31:0] _GEN_4 = 2'h1 == io_INSTR_SEL ? io_rs2 : 32'h0; // @[ZbcExt.scala 100:22 85:18 92:24]
  wire [31:0] _GEN_5 = 2'h1 == io_INSTR_SEL ? CLMULH_io_C_out : _GEN_2; // @[ZbcExt.scala 101:10 92:24]
  wire [31:0] _GEN_6 = 2'h1 == io_INSTR_SEL ? 32'h0 : _GEN_0; // @[ZbcExt.scala 87:18 92:24]
  wire [31:0] _GEN_7 = 2'h1 == io_INSTR_SEL ? 32'h0 : _GEN_1; // @[ZbcExt.scala 88:18 92:24]
  Clmul CLMUL ( // @[ZbcExt.scala 75:21]
    .io_A_in(CLMUL_io_A_in),
    .io_B_in(CLMUL_io_B_in),
    .io_C_out(CLMUL_io_C_out)
  );
  Clmulh CLMULH ( // @[ZbcExt.scala 77:22]
    .io_A_in(CLMULH_io_A_in),
    .io_B_in(CLMULH_io_B_in),
    .io_C_out(CLMULH_io_C_out)
  );
  Clmulr CLMULR ( // @[ZbcExt.scala 79:22]
    .io_A_in(CLMULR_io_A_in),
    .io_B_in(CLMULR_io_B_in),
    .io_C_out(CLMULR_io_C_out)
  );
  assign io_rd = 2'h0 == io_INSTR_SEL ? CLMUL_io_C_out : _GEN_5; // @[ZbcExt.scala 92:24 96:10]
  assign CLMUL_io_A_in = 2'h0 == io_INSTR_SEL ? io_rs1 : 32'h0; // @[ZbcExt.scala 81:17 92:24 94:21]
  assign CLMUL_io_B_in = 2'h0 == io_INSTR_SEL ? io_rs2 : 32'h0; // @[ZbcExt.scala 82:17 92:24 95:21]
  assign CLMULH_io_A_in = 2'h0 == io_INSTR_SEL ? 32'h0 : _GEN_3; // @[ZbcExt.scala 84:18 92:24]
  assign CLMULH_io_B_in = 2'h0 == io_INSTR_SEL ? 32'h0 : _GEN_4; // @[ZbcExt.scala 85:18 92:24]
  assign CLMULR_io_A_in = 2'h0 == io_INSTR_SEL ? 32'h0 : _GEN_6; // @[ZbcExt.scala 87:18 92:24]
  assign CLMULR_io_B_in = 2'h0 == io_INSTR_SEL ? 32'h0 : _GEN_7; // @[ZbcExt.scala 88:18 92:24]
endmodule
